netcdf n20_emissions {
dimensions:
	time = 47;
variables:
        float time(time);
		time:standard_name = "time";
		time:units = "days since 2014-06-06 00:00:00";
	float n2o_control(time);
		n2o_control:long_name = "N2O emissions (control)";
		n2o_control:units = "g N2O-N ha-1 day-1";
		n2o_control:comment = "No standard_name because units are different.";
	float n2o_urea(time);
		n2o_urea:long_name = "N2O emissions (treated with 180 Urea)";
		n2o_urea:units = "g N2O-N ha-1 day-1";
		n2o_urea:comment = "No standard_name because units are different.";
// global attributes:
	:history = "Created on a farm, in the olden days.";
	:Conventions = "CF-1.0";
data:
	time = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46;
	n2o_control = -0.85, 3.25, -0.06, -1.17, 3.59, -2.67, 6.78, -0.42, 0.47, 0.10, -2.33, 2.27, 3.69, -3.89, -2.60, 2.50, 0.79, -2.87, 1.47, 0.75, 2.08, 8.95, -3.24, -4.18, -4.18, 0.20, 4.06, 3.00, 2.34, 2.07, -30.53, -8.87, 30.73, 0.79, 28.68, -1.12, 28.33, 12.25, 2.58, -7.42, 0.44, -1.21, -3.25, -0.47, 3.39, 0.41, -3.06;
	n2o_urea = -0.42, 6.71, 0.34, 4.19, -1.61, -2.36, 5.58, 1.59, -3.53, 1.10, 0.43, 0.39, 5.99, -4.13, -0.24, -2.12, 4.57, -1.93, -0.32, -0.84, 5.48, 3.38, -4.09, 2.45, 2.44, -2.95, -6.11, 8.58, 3.40, -4.16, -6.74, -8.37, 4.91, 0.88, 25.18, -11.32, 21.47, 6.91, 7.86, 4.41, 2.68, -1.39, 0.09, 2.84, 0.98, 0.28, 4.32;
}
